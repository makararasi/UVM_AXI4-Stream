typedef uvm_sequencer #(axi4_seq_item) axi4_seqr;
